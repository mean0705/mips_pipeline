module Shifter( target, shamt, result );
input [31:0] target;
input [4:0] shamt;
output [31:0] result;

wire [31:0] out1, out2, out3, out4;

assign out1[0] = shamt[0] ? 1'b0 : target[0];
assign out1[1] = shamt[0] ? target[0] : target[1];
assign out1[2] = shamt[0] ? target[1] : target[2];
assign out1[3] = shamt[0] ? target[2] : target[3];
assign out1[4] = shamt[0] ? target[3] : target[4];
assign out1[5] = shamt[0] ? target[4] : target[5];
assign out1[6] = shamt[0] ? target[5] : target[6];
assign out1[7] = shamt[0] ? target[6] : target[7];
assign out1[8] = shamt[0] ? target[7] : target[8];
assign out1[9] = shamt[0] ? target[8] : target[9];
assign out1[10] = shamt[0] ? target[9] : target[10];
assign out1[11] = shamt[0] ? target[10] : target[11];
assign out1[12] = shamt[0] ? target[11] : target[12];
assign out1[13] = shamt[0] ? target[12] : target[13];
assign out1[14] = shamt[0] ? target[13] : target[14];
assign out1[15] = shamt[0] ? target[14] : target[15];
assign out1[16] = shamt[0] ? target[15] : target[16];
assign out1[17] = shamt[0] ? target[16] : target[17];
assign out1[18] = shamt[0] ? target[17] : target[18];
assign out1[19] = shamt[0] ? target[18] : target[19];
assign out1[20] = shamt[0] ? target[19] : target[20];
assign out1[21] = shamt[0] ? target[20] : target[21];
assign out1[22] = shamt[0] ? target[21] : target[22];
assign out1[23] = shamt[0] ? target[22] : target[23];
assign out1[24] = shamt[0] ? target[23] : target[24];
assign out1[25] = shamt[0] ? target[24] : target[25];
assign out1[26] = shamt[0] ? target[25] : target[26];
assign out1[27] = shamt[0] ? target[26] : target[27];
assign out1[28] = shamt[0] ? target[27] : target[28];
assign out1[29] = shamt[0] ? target[28] : target[29];
assign out1[30] = shamt[0] ? target[29] : target[30];
assign out1[31] = shamt[0] ? target[30] : target[31];

assign out2[0] = shamt[1] ? 1'b0 : out1[0];
assign out2[1] = shamt[1] ? 1'b0 : out1[1];
assign out2[2] = shamt[1] ? out1[0] : out1[2];
assign out2[3] = shamt[1] ? out1[1] : out1[3];
assign out2[4] = shamt[1] ? out1[2] : out1[4];
assign out2[5] = shamt[1] ? out1[3] : out1[5];
assign out2[6] = shamt[1] ? out1[4] : out1[6];
assign out2[7] = shamt[1] ? out1[5] : out1[7];
assign out2[8] = shamt[1] ? out1[6] : out1[8];
assign out2[9] = shamt[1] ? out1[7] : out1[9];
assign out2[10] = shamt[1] ? out1[8] : out1[10];
assign out2[11] = shamt[1] ? out1[9] : out1[11];
assign out2[12] = shamt[1] ? out1[10] : out1[12];
assign out2[13] = shamt[1] ? out1[11] : out1[13];
assign out2[14] = shamt[1] ? out1[12] : out1[14];
assign out2[15] = shamt[1] ? out1[13] : out1[15];
assign out2[16] = shamt[1] ? out1[14] : out1[16];
assign out2[17] = shamt[1] ? out1[15] : out1[17];
assign out2[18] = shamt[1] ? out1[16] : out1[18];
assign out2[19] = shamt[1] ? out1[17] : out1[19];
assign out2[20] = shamt[1] ? out1[18] : out1[20];
assign out2[21] = shamt[1] ? out1[19] : out1[21];
assign out2[22] = shamt[1] ? out1[20] : out1[22];
assign out2[23] = shamt[1] ? out1[21] : out1[23];
assign out2[24] = shamt[1] ? out1[22] : out1[24];
assign out2[25] = shamt[1] ? out1[23] : out1[25];
assign out2[26] = shamt[1] ? out1[24] : out1[26];
assign out2[27] = shamt[1] ? out1[25] : out1[27];
assign out2[28] = shamt[1] ? out1[26] : out1[28];
assign out2[29] = shamt[1] ? out1[27] : out1[29];
assign out2[30] = shamt[1] ? out1[28] : out1[30];
assign out2[31] = shamt[1] ? out1[29] : out1[31];

assign out3[0] = shamt[2] ? 1'b0 : out2[0];
assign out3[1] = shamt[2] ? 1'b0 : out2[1];
assign out3[2] = shamt[2] ? 1'b0 : out2[2];
assign out3[3] = shamt[2] ? 1'b0 : out2[3];
assign out3[4] = shamt[2] ? out2[0] : out2[4];
assign out3[5] = shamt[2] ? out2[1] : out2[5];
assign out3[6] = shamt[2] ? out2[2] : out2[6];
assign out3[7] = shamt[2] ? out2[3] : out2[7];
assign out3[8] = shamt[2] ? out2[4] : out2[8];
assign out3[9] = shamt[2] ? out2[5] : out2[9];
assign out3[10] = shamt[2] ? out2[6] : out2[10];
assign out3[11] = shamt[2] ? out2[7] : out2[11];
assign out3[12] = shamt[2] ? out2[8] : out2[12];
assign out3[13] = shamt[2] ? out2[9] : out2[13];
assign out3[14] = shamt[2] ? out2[10] : out2[14];
assign out3[15] = shamt[2] ? out2[11] : out2[15];
assign out3[16] = shamt[2] ? out2[12] : out2[16];
assign out3[17] = shamt[2] ? out2[13] : out2[17];
assign out3[18] = shamt[2] ? out2[14] : out2[18];
assign out3[19] = shamt[2] ? out2[15] : out2[19];
assign out3[20] = shamt[2] ? out2[16] : out2[20];
assign out3[21] = shamt[2] ? out2[17] : out2[21];
assign out3[22] = shamt[2] ? out2[18] : out2[22];
assign out3[23] = shamt[2] ? out2[19] : out2[23];
assign out3[24] = shamt[2] ? out2[20] : out2[24];
assign out3[25] = shamt[2] ? out2[21] : out2[25];
assign out3[26] = shamt[2] ? out2[22] : out2[26];
assign out3[27] = shamt[2] ? out2[23] : out2[27];
assign out3[28] = shamt[2] ? out2[24] : out2[28];
assign out3[29] = shamt[2] ? out2[25] : out2[29];
assign out3[30] = shamt[2] ? out2[26] : out2[30];
assign out3[31] = shamt[2] ? out2[27] : out2[31];

assign out4[0] = shamt[3] ? 1'b0 : out3[0];
assign out4[1] = shamt[3] ? 1'b0 : out3[1];
assign out4[2] = shamt[3] ? 1'b0 : out3[2];
assign out4[3] = shamt[3] ? 1'b0 : out3[3];
assign out4[4] = shamt[3] ? 1'b0 : out3[4];
assign out4[5] = shamt[3] ? 1'b0 : out3[5];
assign out4[6] = shamt[3] ? 1'b0 : out3[6];
assign out4[7] = shamt[3] ? 1'b0 : out3[7];
assign out4[8] = shamt[3] ? out3[0] : out3[8];
assign out4[9] = shamt[3] ? out3[1] : out3[9];
assign out4[10] = shamt[3] ? out3[2] : out3[10];
assign out4[11] = shamt[3] ? out3[3] : out3[11];
assign out4[12] = shamt[3] ? out3[4] : out3[12];
assign out4[13] = shamt[3] ? out3[5] : out3[13];
assign out4[14] = shamt[3] ? out3[6] : out3[14];
assign out4[15] = shamt[3] ? out3[7] : out3[15];
assign out4[16] = shamt[3] ? out3[8] : out3[16];
assign out4[17] = shamt[3] ? out3[9] : out3[17];
assign out4[18] = shamt[3] ? out3[10] : out3[18];
assign out4[19] = shamt[3] ? out3[11] : out3[19];
assign out4[20] = shamt[3] ? out3[12] : out3[20];
assign out4[21] = shamt[3] ? out3[13] : out3[21];
assign out4[22] = shamt[3] ? out3[14] : out3[22];
assign out4[23] = shamt[3] ? out3[15] : out3[23];
assign out4[24] = shamt[3] ? out3[16] : out3[24];
assign out4[25] = shamt[3] ? out3[17] : out3[25];
assign out4[26] = shamt[3] ? out3[18] : out3[26];
assign out4[27] = shamt[3] ? out3[19] : out3[27];
assign out4[28] = shamt[3] ? out3[20] : out3[28];
assign out4[29] = shamt[3] ? out3[21] : out3[29];
assign out4[30] = shamt[3] ? out3[22] : out3[30];
assign out4[31] = shamt[3] ? out3[23] : out3[31];

assign result[0] = shamt[4] ? 1'b0 : out4[0];
assign result[1] = shamt[4] ? 1'b0 : out4[1];
assign result[2] = shamt[4] ? 1'b0 : out4[2];
assign result[3] = shamt[4] ? 1'b0 : out4[3];
assign result[4] = shamt[4] ? 1'b0 : out4[4];
assign result[5] = shamt[4] ? 1'b0 : out4[5];
assign result[6] = shamt[4] ? 1'b0 : out4[6];
assign result[7] = shamt[4] ? 1'b0 : out4[7];
assign result[8] = shamt[4] ? 1'b0 : out4[8];
assign result[9] = shamt[4] ? 1'b0 : out4[9];
assign result[10] = shamt[4] ? 1'b0 : out4[10];
assign result[11] = shamt[4] ? 1'b0 : out4[11];
assign result[12] = shamt[4] ? 1'b0 : out4[12];
assign result[13] = shamt[4] ? 1'b0 : out4[13];
assign result[14] = shamt[4] ? 1'b0 : out4[14];
assign result[15] = shamt[4] ? 1'b0 : out4[15];
assign result[16] = shamt[4] ? out4[0] : out4[16];
assign result[17] = shamt[4] ? out4[1] : out4[17];
assign result[18] = shamt[4] ? out4[2] : out4[18];
assign result[19] = shamt[4] ? out4[3] : out4[19];
assign result[20] = shamt[4] ? out4[4] : out4[20];
assign result[21] = shamt[4] ? out4[5] : out4[21];
assign result[22] = shamt[4] ? out4[6] : out4[22];
assign result[23] = shamt[4] ? out4[7] : out4[23];
assign result[24] = shamt[4] ? out4[8] : out4[24];
assign result[25] = shamt[4] ? out4[9] : out4[25];
assign result[26] = shamt[4] ? out4[10] : out4[26];
assign result[27] = shamt[4] ? out4[11] : out4[27];
assign result[28] = shamt[4] ? out4[12] : out4[28];
assign result[29] = shamt[4] ? out4[13] : out4[29];
assign result[30] = shamt[4] ? out4[14] : out4[30];
assign result[31] = shamt[4] ? out4[15] : out4[31];

endmodule